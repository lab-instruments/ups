// -----------------------------------------------------------------------------
//  File Name   :  ups_por.sv
//  Autoher     :  Mike DeLong
//  Date        :  03.16.2019
//  Description :  UPS Power on Reset
// -----------------------------------------------------------------------------
module ups_por(
    // -------------------------------------------------------------------------
    //  Clocks
    // -------------------------------------------------------------------------
    input          clk,

    // -------------------------------------------------------------------------
    //  Clocks
    // -------------------------------------------------------------------------
    input          mode_change,

    // -------------------------------------------------------------------------
    //  Resets
    // -------------------------------------------------------------------------
    output         por_n,
    output         ext_rst_n

);

    // -------------------------------------------------------------------------
    //  Typedefs
    // -------------------------------------------------------------------------
    // -------------------------------------------------------------------------
    //  Variables
    // -------------------------------------------------------------------------
    // State Variable
    logic         por_n_l              = 1'b1;
    logic         ext_rst_n_l          = 1'b1;
    logic [ 7:0]  por_cnt_l            = 8'h0;
    logic [ 7:0]  ext_cnt_l            = 8'h0;

    // -------------------------------------------------------------------------
    //  Pin Assignment Statements
    // -------------------------------------------------------------------------
    assign por_n                       = por_n_l;                               // Power on Reset Assign
    assign ext_rst_n                   = por_n_l & ext_rst_n_l;                 // External Reset Assign

    // -------------------------------------------------------------------------
    //  Generate POR
    // -------------------------------------------------------------------------
    always @(posedge clk) begin : POR_GENERATOR
        if(por_cnt_l < 8'hFF) begin
            por_cnt_l                  <= por_cnt_l + 1'b1;
            por_n_l                    <= 1'b0;

        end else begin
            por_n_l                    <= 1'b1;

        end
    end

    // -------------------------------------------------------------------------
    //  Generate External Reset
    // -------------------------------------------------------------------------
    always @(posedge clk) begin : EXT_RST_GENERATOR
        if (mode_change == 1'b1) begin
            ext_cnt_l                  <= 8'h0;
            ext_rst_n_l                <= 1'b0;

        end else if (ext_cnt_l < 8'hFF) begin
            ext_cnt_l                  <= ext_cnt_l + 1'b1;
            ext_rst_n_l                <= 1'b0;

        end else begin
            ext_rst_n_l                <= 1'b1;

        end
    end

endmodule
