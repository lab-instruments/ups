// -----------------------------------------------------------------------------
//  File Name   :  ups_por.sv
//  Autoher     :  Mike DeLong
//  Date        :  03.16.2019
//  Description :  UPS Power on Reset
// -----------------------------------------------------------------------------
module ups_por(
    // -------------------------------------------------------------------------
    //  Clocks
    // -------------------------------------------------------------------------
    input          clk,

    // -------------------------------------------------------------------------
    //  Power on Reset
    // -------------------------------------------------------------------------
    output         por_n

);

    // -------------------------------------------------------------------------
    //  Typedefs
    // -------------------------------------------------------------------------
    // -------------------------------------------------------------------------
    //  Variables
    // -------------------------------------------------------------------------
    // State Variable
    logic         por_n_l              = 1'b1;
    logic [ 7:0]  por_cnt_l            = 'b0;

    // -------------------------------------------------------------------------
    //  Pin Assignment Statements
    // -------------------------------------------------------------------------
    assign por_n                       = por_n_l;                               // Power on Reset Assign

    // -------------------------------------------------------------------------
    //  Generate POR
    // -------------------------------------------------------------------------
    always @(posedge clk) begin : POR_GENERATOR
        if(por_cnt_l < 8'hFF) begin
            por_cnt_l                  <= por_cnt_l + 1'b1;
            por_n_l                    <= 1'b0;

        end else begin
            por_n_l                    <= 1'b1;

        end
    end

endmodule
